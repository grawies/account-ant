noID	=	"####"
alphabet	=	"abcdefghijklmnopqrstuvwxyzåäöABCDEFGHIJKLMNOPQRSTUVWXYZÅÄÖ"
digits	=	"0123456789"
specialLetters	=	"<>|,;.:-_'*~¨^´`+\?@£$€¥{[]}!"#¤%&/()=µn”“©»«ªßðđŋħłøæ¨þœ→↓←þ®€ł@"
viewMainTitle	=	"Bokföring"
viewMainLoadFilename	=	"Skriv in bokföringsfilens sökväg"
viewMainMenubarEdit	=	"Nytt"
viewMainMenubarEditNewVerificate	=	"Ny verifikation"
viewMainMenubarEditNewVerificateToolTip	=	"Skapa ny verifikation"
viewMainMenubarEditEditVerificate	=	"Visa/Ändra verifikation"
viewMainMenubarEditEditVerificateToolTip	=	"Visa och eventuellt ändra existerande verifikation"
viewMainMenubarViewViewAccount	=	"Visa verifikationer för konto"
viewMainMenubarViewViewAccountToolTip	=	"Visa valt kontos verifikationer"
viewMainMenubarViewToggleActiveAccount	=	"Aktivera/Avaktivera konto"
viewMainMenubarViewToggleActiveAccountToolTip	=	"Ändra kontots status som aktivt eller inaktivt"
viewMainMenubarViewViewEveryAccount	=	"Visa alla konton"
viewMainMenubarViewViewEveryAccountToolTip	=	"Visar både aktiva och inaktiva konton i kontolistan"
viewMainMenubarViewViewActiveAccount	=	"Visa aktiva konton"
viewMainMenubarViewViewActiveAccountToolTip	=	"Visar endast aktiva konton i kontolistan"
viewMainMenubarBudgetNewBudget	=	"Visa budget"
viewMainMenubarBudgetNewBudgetToolTip	=	"Visa/Ändra budgeten för räkenskapsåret"

viewMainAccountplanTabName	=	"Kontoplan"
viewMainVerificatesTabName	=	"Verifikationer"

viewVerificateAccountNum	=	"Konto #"
viewVerificateAccountName	=	"Konto"
viewVerificateDebet	=	"DEBET"
viewVerificateCredit	=	"KREDIT"
viewVerificateChangeSignature	=	"Signatur"
viewVerificateChangeDate	=	"Tidpunkt"
viewVerificateEndOfMonthDescription = "månadsbokslut"

viewVerificateNum	=	"Verifikation #"
viewVerificateDescr	=	"Beskrivning"
viewSum	=	"Summa"
viewVerificateBalance	=	"Balans"

viewVerificateSave	=	"Spara verifikation"
viewBudgetSave	=	"Spara budget"
viewCancel	=	"Stäng"

account	=	"Konto"
viewAccountNum	=	"Kontonummer"
viewAccountVerificate	=	"Visa verifikation"
viewAccountDescription	=	"Kontonamn"
viewBudgetEditMonth	=	"Visa/Ändra månadsbudget"
viewAccountBudget	=	"Visa kontobudget"
editAccountBudget	=	"Månadsfördelning"

viewBudgetTitle	=	"Budget"
viewBudgetMonthDescription	=	"Månad"
viewBudgetMonthBalance	=	"Balans"

report = "Rapport"
viewReportResultsTitle	=	"Resultatrapport"
viewReportBalanceTitle	=	"Balansrapport"
viewMainMenubarReportResultsReport	=	"Resultatrapport"
viewMainMenubarReportResultsReportToolTip	="Generera resultatrapport"
viewMainMenubarReportBalanceReport	=	"Balansrapport"
viewMainMenubarReportBalanceReportToopTip	="Generera balansrapport"
viewSpreadSheetAccountNameEmpty	=	"- - - - - -"

warningVerificateUnbalanced	=	"Obalanserad verifikation"
warningVerificateEmpty	=	"Tomt verifikat"
warningVerificateEmptyText	=	"Inga transaktioner registrerade, verifikationen sparas ej."
warningAmbiguousTransaction	=	"Tvetydig transaktion"
warningAmbiguousTransactionText	=	"En transaktion är otydligt formatterad.
Se till att kontonumret går till ett giltigt konto,
endast en av debet och kredit är ifylld
och eventuell signatur och datum korrekt ifyllda.
Alternativt se till att raden är tom.
Gäller rad "
warningNewVerificateAlreadyOpen	=	"Avsluta pågående ny verifikation"
warningNewVerificateAlreadyOpenText	=	"En fönster för ny verifikation är redan öppet.
Avsluta det nuvarande om du vill öppna ett nytt."

period = "Period:"
forPeriod = " för perioden "
columns = "Kolumner:"
date = "Datum:"
warningWrongFormatDateTitle = "Ogiltigt datum"
warningWrongFormatDate	=	"Felformaterat datum, skall vara på formen YYYY-MM-DD"
warningWrongFormatDateFiscal = " och ligga inom verksamhetsåret."
warningLoadFileNotFound	=	"Ogiltig sökväg!"
warningLoadFileNotFoundText	=	"Filens sökväg hittades inte"

showSpecificAccounts = "Visa kontospecifikation"

warningbudgetWindowAlreadyOpen	=	"Nytt budgetfönster kan ej öppnas"
warningbudgetWindowAlreadyOpenText	=	"Budgeten syns och används redan i ett annat fönster."
save	=	"Spara"
saveToolTip	=	"Spara fil till disk"
load	=	"Öppna"
loadToolTip	=	"Ladda in en fil från disk"
exit	=	"Avsluta"
exitToolTip	=	"Avsluta programmet utan att spara"
viewMonth0	=	"januari"
viewMonth1	=	"februari"
viewMonth2	=	"mars"
viewMonth3	=	"april"
viewMonth4	=	"maj"
viewMonth5	=	"juni"
viewMonth6	=	"juli"
viewMonth7	=	"augusti"
viewMonth8	=	"september"
viewMonth9	=	"oktober"
viewMonth10	=	"november"
viewMonth11	=	"december"

showReportInWindow = "Bildskärm"
showReportInBrowser = "Webbläsare"
saveReportAsHTML = "Spara HTML..."
saveReportAsPDF = "Spara PDF..."
sendReportToPrinter = "Utskrift..."

showPeriodColumn = "Period"
showAccumulatedColumn = "Ackumulerat"
showLastYearColumn = "Föregående år"
showBudgetColumn = "Budget"
showPeriodBudgetQuotientColumn = "Visa period/budget"

showBudget = "Budget"
showLastYear = "Föregående år"
showWholeYears = "Helår"
showAccumulated = "Ackumulerat"
showPeriod = "Period"

preliminary = "Preliminär"

saveBeforeExit = "Vill du spara innan du avslutar?"
saveBeforeExitTitle = "Avsluta program"

resultReportSubTitlePreliminary = "Preliminär"
resultReportColumnTitleAccountID = "Konto #"
resultReportColumnTitleAccountName = "Kontonamn"
resultReportColumnTitlePeriod = "Period"
resultReportColumnTitleAccumulated = "Ackumulerat"
resultReportColumnTitleLastYearPeriod = "Fjolår period"
resultReportColumnTitleLastYearAccumulated = "Fjolår ackumulerat"
resultReportColumnTitleLastYearFiscalYear = "Fjolår räkenskapsår"
resultReportColumnTitleBudgetPeriod = "Budget period"
resultReportColumnTitleBudgetAccumulated = "Budget ackumulerat"
resultReportColumnTitleBudgetFiscalYear = "Budget räkenskapsår"
resultReportColumnTitlePeriodBudgetQuotient = "Period/budget"

accountPlan_1 = "Tillgångar"
accountPlan_10 = "Immateriella anläggningstillgångar"
accountPlan_11 = "Byggnader och mark"
accountPlan_12 = "Maskiner och inventarier"
accountPlan_13 = "Finansiella anläggningstillgångar"
accountPlan_14 = "Lager, produkter i arbete och pågpende arbeten"
accountPlan_15 = "Kundfordringar"
accountPlan_16 = "Övriga kortfristiga fordringar"
accountPlan_17 = "Förutbetalda kostnader och upplupna intäkter"
accountPlan_18 = "Kortfristiga placeringar"
accountPlan_19 = "Kassa och bank"
accountPlan_2 = "Eget kapital, avsättningar och skulder"
accountPlan_20 = "Eget kapital"
accountPlan_21 = "Obeskattade reserver"
accountPlan_22 = "Avsättningar"
accountPlan_23 = "Långfristiga skulder"
accountPlan_24 = "Kortfristiga skulder till kreditinstitut, kunder och leverantörer"
accountPlan_25 = "Skatteskulder"
accountPlan_26 = "Moms och särskilda punktskatter"
accountPlan_27 = "Personalens skatter, avgifter och löneavdrag"
accountPlan_28 = "Övriga kortfristiga skulder"
accountPlan_29 = "Upplupna kostnader och förutbetalda intäkter"
accountPlan_3 = "Rörelsens inkomster/intäkter"
accountPlan_30 = "Huvudintäkter"
accountPlan_31 = "Huvudintäkter"
accountPlan_32 = "Huvudintäkter"
accountPlan_34 = "Huvudintäkter"
accountPlan_35 = "Fakturerade kostnader"
accountPlan_36 = "Rörelsens sidointäkter"
accountPlan_37 = "Intäktskorrigeringar"
accountPlan_38 = "Aktiverat arbete för egen räkning"
accountPlan_39 = "Övriga rörelseintäkter"
accountPlan_4 = "Utgifter/kostnader för varor, material och vissa köpta tjänster"
accountPlan_40 = "Inköp av varor och material"
accountPlan_41 = "Inköp av varor och material"
accountPlan_42 = "Inköp av varor och material"
accountPlan_43 = "Inköp av varor och material"
accountPlan_44 = "Inköp av varor och material"
accountPlan_45 = "Inköp av varor och material"
accountPlan_46 = "Legoarbeten, underentreprenader"
accountPlan_47 = "Reduktion av inköpspriser"
accountPlan_48 = "(Fri kontogrupp)"
accountPlan_49 = "Förändrigar av lager, produkter i arbeten och pågående arbeten"
accountPlan_5 = "Övriga externa rörelseutgifter/kostnader"
accountPlan_50 = "Lokalkostnader"
accountPlan_51 = "Fastighetskostnader"
accountPlan_52 = "Hyra av anälggningstillgångar"
accountPlan_53 = "Energikostnader"
accountPlan_54 = "Förbrukningsinventarier och förbrukningsmaterial"
accountPlan_55 = "Reparation och underhåll"
accountPlan_56 = "Kostnader för transportmedel"
accountPlan_57 = "Frakter och transporter"
accountPlan_58 = "Resekostnader"
accountPlan_59 = "Reklam och PR"
accountPlan_6 = "Övriga externa rörelseutgifter/kostnader"
accountPlan_60 = "Övriga försäljningskostnader"
accountPlan_61 = "Kontorsmateriel och trycksaker"
accountPlan_62 = "Tele och post"
accountPlan_63 = "Företagsförsäkringar och övriga riskkostnader"
accountPlan_64 = "Förvaltningskostnader"
accountPlan_65 = "Övriga externa tjänster"
accountPlan_66 = "(Fri kontogrupp)"
accountPlan_67 = "(Fri kontogrupp)"
accountPlan_68 = "Inhyrd personal"
accountPlan_69 = "Övriga externa kostnader"
accountPlan_7 = "Utgifter/kostnader för personal, avskrivningar m.m."
accountPlan_70 = "Löner till kollektivanställda"
accountPlan_71 = "(Fri kontogrupp)"
accountPlan_72 = "Löner till tjänstemän och företagsledare"
accountPlan_73 = "Kostnadsersättningar och förmåner"
accountPlan_74 = "Pensionskostnader"
accountPlan_75 = "Sociala och andra avgifter enligt lag och avtal"
accountPlan_76 = "Övriga personalkostnader"
accountPlan_77 = "Nedskrivningar och återföring av nedskrivningar"
accountPlan_78 = "Avskrivningar enligt plan"
accountPlan_79 = "Övriga rörelsekostnader"
accountPlan_8 = "Finansiella och andra inkomster/intäkter och utgifter/kostnader"
accountPlan_80 = "Resultat från andelar i koncernföretag"
accountPlan_81 = "Resultat från andelar i intresseföretag"
accountPlan_82 = "Resultat från övriga värdepapper och långfristiga fordringar (anläggningstillgångar)"
accountPlan_83 = "Övriga ränkteintäkter och liknande resultatposter"
accountPlan_84 = "Räntekostnader och liknande resultatposter"
accountPlan_85 = "(Fri kontogrupp)"
accountPlan_86 = "(Fri kontogrupp)"
accountPlan_87 = "Extraordinära intäkter och kostnader"
accountPlan_88 = "Bokslutsdispositioner"
accountPlan_89 = "Skatter och årets resultat"

